module accumulator(
  input        clk, reset, req, 
  output logic done);