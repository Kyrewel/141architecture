// cache memory/register file
// default address pointer width = 4, for 16 registers
module reg_file #(parameter pw=4)(
  input[7:0] dat_in,
  input      clk,
  input      wr_en,           // write enable
  input[pw-1:0] wr_addr,		  // write address pointer
              rd_addrA,		  // read address pointers
			  rd_addrB,
  input wire [11:0] prog_ctr,
  output logic[7:0] datA_out, // read data
                    datB_out);
					
  logic [11:0] oldPC = -1;

  logic [7:0] core[2**pw];    // 2-dim array  8 wide  16 deep

// reads are combinational
  assign datA_out = core[rd_addrA];
  assign datB_out = core[rd_addrB];

// writes are sequential (clocked)
  always_ff @(posedge clk) begin
    if(wr_en && oldPC !== prog_ctr) begin				   // anything but stores or no ops
      $display("RF: time=%t writing %d to reg %d", $time, dat_in, wr_addr); 
      core[wr_addr] <= dat_in;
	    oldPC <= prog_ctr;
	  end	
  end
  // Debugging code to print the contents of the core register array
  logic [7:0] old_core[2**pw]; // Array to store old values of core for comparison

  initial begin
    for (int i = 0; i < 2**pw; i++) begin
      old_core[i] = 'bx; // Initialize old_core values
    end
  end

  always_ff @(posedge clk) begin
    for (int i = 0; i < 2**pw; i++) begin
      if (core[i] !== old_core[i]) begin
        $display("RF: core[%0d] changed to %d at time %t", i, core[i], $time);
        for (int j = 0; j < 2**pw; j++) begin
          $display("RF: core[%0d] = %d", j, core[j]);
        end
        old_core = core; // Update old_core to the current state
        break;
      end
    end
  end

endmodule
/*
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
	  xxxx_xxxx
*/