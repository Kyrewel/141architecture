put 0       0000 0000 1
put 1       0000 0001 1
ld          0000 0001 1


put 1       0000 0001 1
put 1       0000 0001 1
ld          0000 0001 0

put 2       0000 0010 1
put 0       0000 0000 1
put 1       0000 0001 1

add         0000 1010 0