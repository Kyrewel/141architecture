put 0
put 1    
ld


put 1
put 1
ld

put 2
put 0
put 1

add